.title KiCad schematic
.model __M8 NMOS level=8
.model __M12 NMOS level=8
.model __M9 NMOS level=8
.model __M5 NMOS level=8
.model __M11 NMOS level=8
.model __M10 NMOS level=8
.model __M6 NMOS level=8
.model __M7 NMOS level=8
.model __M4 PMOS level=8
.model __M2 PMOS level=8
.model __M1 PMOS level=8
.model __M3 PMOS level=8
M8 Net-_M4-D_ Net-_M6-B_ Net-_M12-D_ Net-_M12-D_ __M8
M12 Net-_M12-D_ Net-_M11-D_ eSim_GND eSim_GND __M12
M9 Net-_M10-G_ Net-_M10-G_ eSim_GND eSim_GND __M9
M5 Iin Iin Net-_M10-G_ Net-_M10-G_ __M5
R2 Iout_RG Iout 330
M11 Net-_M11-D_ Net-_M10-B_ eSim_GND eSim_GND __M11
M10 Net-_M10-D_ Net-_M10-G_ eSim_GND Net-_M10-B_ __M10
M6 Net-_M3-D_ Iin Net-_M10-D_ Net-_M6-B_ __M6
M7 Iout Net-_M4-D_ Net-_M11-D_ Net-_M11-D_ __M7
M4 Net-_M4-D_ Net-_M3-D_ Net-_M2-D_ Net-_M2-D_ __M4
M2 Net-_M2-D_ Net-_M1-D_ eSim_VCC eSim_VCC __M2
R1 Iin Iin_r 330
M1 Net-_M1-D_ Net-_M1-D_ eSim_VCC eSim_VCC __M1
Vv1 Iin_r Iout_RG DC 4 
M3 Net-_M3-D_ Net-_M3-D_ Net-_M1-D_ Net-_M1-D_ __M3
.end
